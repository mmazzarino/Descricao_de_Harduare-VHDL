----------------------------------------------------------------------------------
-- Course: Engenharia de Controle e Automa��o
-- Subject: Laborat�rio de Circu�tos L�gicos II
-- Engineer: Matheus Mazzarino
-- Create Date: Outubro 2018 
-- Module Name: DISPLAY_LCD_16X2 - ARQ_DISPLAY_LCD_16X2 

-- Description: 

----------------------------------------------------------------------------------
library IEEE;
library UNISIM;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_ARITH.ALL; 
use UNISIM.VComponents.all;

entity DISPLAY_LCD_16X2 is
end DISPLAY_LCD_16X2;

architecture ARQ_DISPLAY_LCD_16X2 of DISPLAY_LCD_16X2 is

begin


end ARQ_DISPLAY_LCD_16X2;

